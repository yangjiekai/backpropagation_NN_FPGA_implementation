library verilog;
use verilog.vl_types.all;
entity TopTest is
end TopTest;
